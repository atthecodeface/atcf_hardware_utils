/** @copyright (C) 2020,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   fifo_status.cdl
 * @brief  A FIFO status recording module
 *
 */
/*a Constants */
constant integer fifo_depth_max=16;
constant integer fifo_entries_mask=(1<<sizeof(fifo_depth_max))-1;

include "fifo_status.h"

/*a Module
 */
module fifo_status( clock clk                            "Clock for logic",
                    input bit reset_n                    "Active low reset",
                    input bit push,
                    input bit pop,
                    input bit[32] max_entries "Should be hardwired in parent",
                    output t_fifo_status fifo_status
    )
{
    /*b State etc  */
    default reset active_low reset_n;
    default clock clk;

    clocked t_fifo_status fifo_status={*=0, empty=1}  "Fifo status";

    /*b Status logic */
    status_logic """
    """: {
        fifo_status.pushed <= push;
        fifo_status.popped <= pop;
        if (fifo_status.empty && pop && !push) {
            assert(0, "Fifo underflowed");
            fifo_status.underflowed <= 1;
        }
        if (fifo_status.full && push && !pop) {
            assert(0, "Fifo overflowed");
            fifo_status.overflowed <= 1;
        }
        if (pop) {
            if (push) {
                fifo_status.entries_full <= fifo_status.entries_full & fifo_entries_mask;
            } else {
                fifo_status.full <= 0;
                fifo_status.entries_full <= (fifo_status.entries_full-1) & fifo_entries_mask;
                if (fifo_status.entries_full==1) {
                    fifo_status.empty <= 1;
                }
            }
        } else {
            if (push) {
                fifo_status.empty <= 0;
                fifo_status.entries_full <= (fifo_status.entries_full+1) & fifo_entries_mask;
                if (fifo_status.entries_full==max_entries-1) {
                    fifo_status.full <= 1;
                }
            }
        }
        
        /*b All done */
    }

    /*b All done */
}
