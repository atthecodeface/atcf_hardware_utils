/** Copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *   http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * @file  tb_teletext.cdl
 * @brief Testbench for teletext decoder module
 *
 * This is a simple testbench for the teletext decoder.
 */
/*a Includes */
include "dprintf.h"
include "dprintf_modules.h"

/*a External modules */
extern module se_test_harness( clock clk,
                               output bit[4] reqs,
                               input bit[4] acks,
                               input t_dprintf_byte dprintf_byte
    )
{
    timing from rising clock clk reqs;
    timing to   rising clock clk acks, dprintf_byte;
}

/*a Module */
module tb_dprintf_mux( clock clk,
                       input bit reset_n
)
{

    /*b Nets */
    net bit[4] reqs;
    //net bit[4] acks;
    net t_dprintf_req_2   req_01;
    net t_dprintf_req_2   req_012;
    comb t_dprintf_req_4  req_012b;
    net t_dprintf_req_4   req_0123;
    net bit             ack_0;
    net bit             ack_1;
    net bit             ack_2;
    net bit             ack_3;
    net bit             ack_01;
    net bit             ack_012;
    net bit             ack_0123;
    net t_dprintf_byte dprintf_byte;
    comb t_dprintf_req_2   req_0;
    comb t_dprintf_req_2   req_1;
    comb t_dprintf_req_2   req_2;
    comb t_dprintf_req_4   req_3;

    /*b Instantiations */
    instantiations: {
        req_0 = {valid=reqs[0], address=0x1010, data_0=64h41_42_43_44_45_46_47_48, data_1=64h_83_de_ad_83_be_ef_ff_00 };
        req_1 = {valid=reqs[1], address=0x2010, data_0=64h20_ff_0000_00000000, data_1=0};
        req_2 = {valid=reqs[2], address=0x3010, data_0=64h22_ff_0000_00000000, data_1=0};
        req_3 = {valid=reqs[3], address=0x4010, data_0=64h33_00_0000_00000000, data_1=0, data_2=64h34_00_0000_00000000, data_3=64h00000000_000000_35};
        se_test_harness th( clk <- clk,
                            reqs => reqs,
                            acks <= bundle(ack_3, ack_2, ack_1, ack_0),
                            dprintf_byte <=  dprintf_byte
                                );
        
        dprintf_2_mux mux01( clk <- clk,
                                   reset_n <= reset_n,
                                   req_a <= req_0,
                                   req_b <= req_1,
                                   ack_a => ack_0,
                                   ack_b => ack_1,
                                   req => req_01,
                                   ack <= ack_01 );

        dprintf_2_mux mux012( clk <- clk,
                                   reset_n <= reset_n,
                                   req_a <= req_01,
                                   req_b <= req_2,
                                   ack_a => ack_01,
                                   ack_b => ack_2,
                                   req => req_012,
                                   ack <= ack_012 );

        req_012b = {valid   = req_012.valid,
                    address = req_012.address,
                    data_0  = req_012.data_0,
                    data_1  = req_012.data_1,
                    data_2  = -1,
                    data_3  = -1};
                    
        dprintf_4_mux mux013( clk <- clk,
                                   reset_n <= reset_n,
                                   req_a <= req_012b,
                                   req_b <= req_3,
                                   ack_a => ack_012,
                                   ack_b => ack_3,
                                   req => req_0123,
                                   ack <= ack_0123 );

        dprintf dut( clk <- clk,
                              reset_n <= reset_n,
                              dprintf_req <= req_0123,
                              dprintf_ack => ack_0123,
                              dprintf_byte =>  dprintf_byte
            );
    }

    /*b All done */
}
